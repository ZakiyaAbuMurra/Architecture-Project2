module CPU(clk, inst_Din);
	input clk;
	input [31:0] inst_Din;
	
	wire [31:0] next_pc0, next_pc1, next_pc2; 
	
	
	
	
	
	
endmodule