`include "sign_extender.v"
`include "stack.v"
`include "mux_2x1.v"
`include "RegFile.v"
`include "mux4x1.v"
`include "InstMem.v"
`include "IR.v"
`include "DataMem.v"
`include "ControlUnit.v"
`include  "ALU.v"
`include "pc.v"
`include "dff.v"
`include "adder.v"
`include "cpu.v"

